module group_detection (
    input iColor,
    input iDVAL,
    input iX_Cont,
    input iY_Cont,
    output oX,
    output oY,
    output oDVAL,
    input iCLK,
    input iRST
);


endmodule