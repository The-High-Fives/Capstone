module IPU();

endmodule