module cpu
(
    input clk,
    input rst_n
);

endmodule